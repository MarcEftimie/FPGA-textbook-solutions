module time_multiplexer(
    input wire clk_i,
    input wire rst_i,
    input wire [7:0] in0, in1, in2, in3,
    output logic [3:0] an,
    output logic [7:0] sseg
);

    // Declarations
endmodule