module dual_priority_encoder(
    
);

endmodule